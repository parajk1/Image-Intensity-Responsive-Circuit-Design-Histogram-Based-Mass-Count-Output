module mux255 # (parameter WIDTH = 8)
(input [WIDTH-1:0] d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,
d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,d33,d34,d35,d36,d37,d38,d39,d40,d41,
d42,d43,d44,d45,d46,d47,d48,d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61,d62,d63,d64,d65,d66,d67,d68,
d69,d70,d71,d72,d73,d74,d75,d76,d77,d78,d79,d80,d81,d82,d83,d84,d85,d86,d87,d88,d89,d90,d91,d92,d93,d94,d95,
d96,d97,d98,d99,d100,d101,d102,d103,d104,d105,d106,d107,d108,d109,d110,d111,d112,d113,d114,d115,d116,d117,d118,
d119,d120,d121,d122,d123,d124,d125,d126,d127,d128,d129,d130,d131,d132,d133,d134,d135,d136,d137,d138,d139,d140,d141,
d142,d143,d144,d145,d146,d147,d148,d149,d150,d151,d152,d153,d154,d155,d156,d157,d158,d159,d160,d161,d162,d163,d164,
d165,d166,d167,d168,d169,d170,d171,d172,d173,d174,d175,d176,d177,d178,d179,d180,d181,d182,d183,d184,d185,d186,d187,
d188,d189,d190,d191,d192,d193,d194,d195,d196,d197,d198,d199,d200,d201,d202,d203,d204,d205,d206,d207,d208,d209,d210,
d211,d212,d213,d214,d215,d216,d217,d218,d219,d220,d221,d222,d223,d224,d225,d226,d227,d228,d229,d230,d231,d232,d233,
d234,d235,d236,d237,d238,d239,d240,d241,d242,d243,d244,d245,d246,d247,d248,d249,d250,d251,d252,d253,d254,d255,
input[7:0] s,
output reg [WIDTH-1:0] y);
always @ (*) begin

case(s)
8'b00000000 : y = d0;
8'b00000001 : y = d1;
8'b00000010 : y = d2;
8'b00000011 : y = d3;
8'b00000100 : y = d4;
8'b00000101 : y = d5;
8'b00000110 : y = d6;
8'b00000111 : y = d7;
8'b00001000 : y = d8;
8'b00001001 : y = d9;
8'b00001010 : y = d10;
8'b00001011 : y = d11;
8'b00001100 : y = d12;
8'b00001101 : y = d13;
8'b00001110 : y = d14;
8'b00001111 : y = d15;
8'b00010000 : y = d16;
8'b00010001 : y = d17;
8'b00010010 : y = d18;
8'b00010011 : y = d19;
8'b00010100 : y = d20;
8'b00010101 : y = d21;
8'b00010110 : y = d22;
8'b00010111 : y = d23;
8'b00011000 : y = d24;
8'b00011001 : y = d25;
8'b00011010 : y = d26;
8'b00011011 : y = d27;
8'b00011100 : y = d28;
8'b00011101 : y = d29;
8'b00011110 : y = d30;
8'b00011111 : y = d31;
8'b00100000 : y = d32;
8'b00100001 : y = d33;
8'b00100010 : y = d34;
8'b00100011 : y = d35;
8'b00100100 : y = d36;
8'b00100101 : y = d37;
8'b00100110 : y = d38;
8'b00100111 : y = d39;
8'b00101000 : y = d40;
8'b00101001 : y = d41;
8'b00101010 : y = d42;
8'b00101011 : y = d43;
8'b00101100 : y = d44;
8'b00101101 : y = d45;
8'b00101110 : y = d46;
8'b00101111 : y = d47;
8'b00110000 : y = d48;
8'b00110001 : y = d49;
8'b00110010 : y = d50;
8'b00110011 : y = d51;
8'b00110100 : y = d52;
8'b00110101 : y = d53;
8'b00110110 : y = d54;
8'b00110111 : y = d55;
8'b00111000 : y = d56;
8'b00111001 : y = d57;
8'b00111010 : y = d58;
8'b00111011 : y = d59;
8'b00111100 : y = d60;
8'b00111101 : y = d61;
8'b00111110 : y = d62;
8'b00111111 : y = d63;
8'b01000000 : y = d64;
8'b01000001 : y = d65;
8'b01000010 : y = d66;
8'b01000011 : y = d67;
8'b01000100 : y = d68;
8'b01000101 : y = d69;
8'b01000110 : y = d70;
8'b01000111 : y = d71;
8'b01001000 : y = d72;
8'b01001001 : y = d73;
8'b01001010 : y = d74;
8'b01001011 : y = d75;
8'b01001100 : y = d76;
8'b01001101 : y = d77;
8'b01001110 : y = d78;
8'b01001111 : y = d79;
8'b01010000 : y = d80;
8'b01010001 : y = d81;
8'b01010010 : y = d82;
8'b01010011 : y = d83;
8'b01010100 : y = d84;
8'b01010101 : y = d85;
8'b01010110 : y = d86;
8'b01010111 : y = d87;
8'b01011000 : y = d88;
8'b01011001 : y = d89;
8'b01011010 : y = d90;
8'b01011011 : y = d91;
8'b01011100 : y = d92;
8'b01011101 : y = d93;
8'b01011110 : y = d94;
8'b01011111 : y = d95;
8'b01100000 : y = d96;
8'b01100001 : y = d97;
8'b01100010 : y = d98;
8'b01100011 : y = d99;
8'b01100100 : y = d100;
8'b01100101 : y = d101;
8'b01100110 : y = d102;
8'b01100111 : y = d103;
8'b01101000 : y = d104;
8'b01101001 : y = d105;
8'b01101010 : y = d106;
8'b01101011 : y = d107;
8'b01101100 : y = d108;
8'b01101101 : y = d109;
8'b01101110 : y = d110;
8'b01101111 : y = d111;
8'b01110000 : y = d112;
8'b01110001 : y = d113;
8'b01110010 : y = d114;
8'b01110011 : y = d115;
8'b01110100 : y = d116;
8'b01110101 : y = d117;
8'b01110110 : y = d118;
8'b01110111 : y = d119;
8'b01111000 : y = d120;
8'b01111001 : y = d121;
8'b01111010 : y = d122;
8'b01111011 : y = d123;
8'b01111100 : y = d124;
8'b01111101 : y = d125;
8'b01111110 : y = d126;
8'b01111111 : y = d127;
8'b10000000 : y = d128;
8'b10000001 : y = d129;
8'b10000010 : y = d130;
8'b10000011 : y = d131;
8'b10000100 : y = d132;
8'b10000101 : y = d133;
8'b10000110 : y = d134;
8'b10000111 : y = d135;
8'b10001000 : y = d136;
8'b10001001 : y = d137;
8'b10001010 : y = d138;
8'b10001011 : y = d139;
8'b10001100 : y = d140;
8'b10001101 : y = d141;
8'b10001110 : y = d142;
8'b10001111 : y = d143;
8'b10010000 : y = d144;
8'b10010001 : y = d145;
8'b10010010 : y = d146;
8'b10010011 : y = d147;
8'b10010100 : y = d148;
8'b10010101 : y = d149;
8'b10010110 : y = d150;
8'b10010111 : y = d151;
8'b10011000 : y = d152;
8'b10011001 : y = d153;
8'b10011010 : y = d154;
8'b10011011 : y = d155;
8'b10011100 : y = d156;
8'b10011101 : y = d157;
8'b10011110 : y = d158;
8'b10011111 : y = d159;
8'b10100000 : y = d160;
8'b10100001 : y = d161;
8'b10100010 : y = d162;
8'b10100011 : y = d163;
8'b10100100 : y = d164;
8'b10100101 : y = d165;
8'b10100110 : y = d166;
8'b10100111 : y = d167;
8'b10101000 : y = d168;
8'b10101001 : y = d169;
8'b10101010 : y = d170;
8'b10101011 : y = d171;
8'b10101100 : y = d172;
8'b10101101 : y = d173;
8'b10101110 : y = d174;
8'b10101111 : y = d175;
8'b10110000 : y = d176;
8'b10110001 : y = d177;
8'b10110010 : y = d178;
8'b10110011 : y = d179;
8'b10110100 : y = d180;
8'b10110101 : y = d181;
8'b10110110 : y = d182;
8'b10110111 : y = d183;
8'b10111000 : y = d184;
8'b10111001 : y = d185;
8'b10111010 : y = d186;
8'b10111011 : y = d187;
8'b10111100 : y = d188;
8'b10111101 : y = d189;
8'b10111110 : y = d190;
8'b10111111 : y = d191;
8'b11000000 : y = d192;
8'b11000001 : y = d193;
8'b11000010 : y = d194;
8'b11000011 : y = d195;
8'b11000100 : y = d196;
8'b11000101 : y = d197;
8'b11000110 : y = d198;
8'b11000111 : y = d199;
8'b11001000 : y = d200;
8'b11001001 : y = d201;
8'b11001010 : y = d202;
8'b11001011 : y = d203;
8'b11001100 : y = d204;
8'b11001101 : y = d205;
8'b11001110 : y = d206;
8'b11001111 : y = d207;
8'b11010000 : y = d208;
8'b11010001 : y = d209;
8'b11010010 : y = d210;
8'b11010011 : y = d211;
8'b11010100 : y = d212;
8'b11010101 : y = d213;
8'b11010110 : y = d214;
8'b11010111 : y = d215;
8'b11011000 : y = d216;
8'b11011001 : y = d217;
8'b11011010 : y = d218;
8'b11011011 : y = d219;
8'b11011100 : y = d220;
8'b11011101 : y = d221;
8'b11011110 : y = d222;
8'b11011111 : y = d223;
8'b11100000 : y = d224;
8'b11100001 : y = d225;
8'b11100010 : y = d226;
8'b11100011 : y = d227;
8'b11100100 : y = d228;
8'b11100101 : y = d229;
8'b11100110 : y = d230;
8'b11100111 : y = d231;
8'b11101000 : y = d232;
8'b11101001 : y = d233;
8'b11101010 : y = d234;
8'b11101011 : y = d235;
8'b11101100 : y = d236;
8'b11101101 : y = d237;
8'b11101110 : y = d238;
8'b11101111 : y = d239;
8'b11110000 : y = d240;
8'b11110001 : y = d241;
8'b11110010 : y = d242;
8'b11110011 : y = d243;
8'b11110100 : y = d244;
8'b11110101 : y = d245;
8'b11110110 : y = d246;
8'b11110111 : y = d247;
8'b11111000 : y = d248;
8'b11111001 : y = d249;
8'b11111010 : y = d250;
8'b11111011 : y = d251;
8'b11111100 : y = d252;
8'b11111101 : y = d253;
8'b11111110 : y = d254;
8'b11111111 : y = d255;
default : y=256'bx;
endcase
end
endmodule