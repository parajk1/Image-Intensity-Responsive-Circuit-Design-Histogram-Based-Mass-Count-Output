library verilog;
use verilog.vl_types.all;
entity mux255 is
    generic(
        WIDTH           : integer := 8
    );
    port(
        d0              : in     vl_logic_vector;
        d1              : in     vl_logic_vector;
        d2              : in     vl_logic_vector;
        d3              : in     vl_logic_vector;
        d4              : in     vl_logic_vector;
        d5              : in     vl_logic_vector;
        d6              : in     vl_logic_vector;
        d7              : in     vl_logic_vector;
        d8              : in     vl_logic_vector;
        d9              : in     vl_logic_vector;
        d10             : in     vl_logic_vector;
        d11             : in     vl_logic_vector;
        d12             : in     vl_logic_vector;
        d13             : in     vl_logic_vector;
        d14             : in     vl_logic_vector;
        d15             : in     vl_logic_vector;
        d16             : in     vl_logic_vector;
        d17             : in     vl_logic_vector;
        d18             : in     vl_logic_vector;
        d19             : in     vl_logic_vector;
        d20             : in     vl_logic_vector;
        d21             : in     vl_logic_vector;
        d22             : in     vl_logic_vector;
        d23             : in     vl_logic_vector;
        d24             : in     vl_logic_vector;
        d25             : in     vl_logic_vector;
        d26             : in     vl_logic_vector;
        d27             : in     vl_logic_vector;
        d28             : in     vl_logic_vector;
        d29             : in     vl_logic_vector;
        d30             : in     vl_logic_vector;
        d31             : in     vl_logic_vector;
        d32             : in     vl_logic_vector;
        d33             : in     vl_logic_vector;
        d34             : in     vl_logic_vector;
        d35             : in     vl_logic_vector;
        d36             : in     vl_logic_vector;
        d37             : in     vl_logic_vector;
        d38             : in     vl_logic_vector;
        d39             : in     vl_logic_vector;
        d40             : in     vl_logic_vector;
        d41             : in     vl_logic_vector;
        d42             : in     vl_logic_vector;
        d43             : in     vl_logic_vector;
        d44             : in     vl_logic_vector;
        d45             : in     vl_logic_vector;
        d46             : in     vl_logic_vector;
        d47             : in     vl_logic_vector;
        d48             : in     vl_logic_vector;
        d49             : in     vl_logic_vector;
        d50             : in     vl_logic_vector;
        d51             : in     vl_logic_vector;
        d52             : in     vl_logic_vector;
        d53             : in     vl_logic_vector;
        d54             : in     vl_logic_vector;
        d55             : in     vl_logic_vector;
        d56             : in     vl_logic_vector;
        d57             : in     vl_logic_vector;
        d58             : in     vl_logic_vector;
        d59             : in     vl_logic_vector;
        d60             : in     vl_logic_vector;
        d61             : in     vl_logic_vector;
        d62             : in     vl_logic_vector;
        d63             : in     vl_logic_vector;
        d64             : in     vl_logic_vector;
        d65             : in     vl_logic_vector;
        d66             : in     vl_logic_vector;
        d67             : in     vl_logic_vector;
        d68             : in     vl_logic_vector;
        d69             : in     vl_logic_vector;
        d70             : in     vl_logic_vector;
        d71             : in     vl_logic_vector;
        d72             : in     vl_logic_vector;
        d73             : in     vl_logic_vector;
        d74             : in     vl_logic_vector;
        d75             : in     vl_logic_vector;
        d76             : in     vl_logic_vector;
        d77             : in     vl_logic_vector;
        d78             : in     vl_logic_vector;
        d79             : in     vl_logic_vector;
        d80             : in     vl_logic_vector;
        d81             : in     vl_logic_vector;
        d82             : in     vl_logic_vector;
        d83             : in     vl_logic_vector;
        d84             : in     vl_logic_vector;
        d85             : in     vl_logic_vector;
        d86             : in     vl_logic_vector;
        d87             : in     vl_logic_vector;
        d88             : in     vl_logic_vector;
        d89             : in     vl_logic_vector;
        d90             : in     vl_logic_vector;
        d91             : in     vl_logic_vector;
        d92             : in     vl_logic_vector;
        d93             : in     vl_logic_vector;
        d94             : in     vl_logic_vector;
        d95             : in     vl_logic_vector;
        d96             : in     vl_logic_vector;
        d97             : in     vl_logic_vector;
        d98             : in     vl_logic_vector;
        d99             : in     vl_logic_vector;
        d100            : in     vl_logic_vector;
        d101            : in     vl_logic_vector;
        d102            : in     vl_logic_vector;
        d103            : in     vl_logic_vector;
        d104            : in     vl_logic_vector;
        d105            : in     vl_logic_vector;
        d106            : in     vl_logic_vector;
        d107            : in     vl_logic_vector;
        d108            : in     vl_logic_vector;
        d109            : in     vl_logic_vector;
        d110            : in     vl_logic_vector;
        d111            : in     vl_logic_vector;
        d112            : in     vl_logic_vector;
        d113            : in     vl_logic_vector;
        d114            : in     vl_logic_vector;
        d115            : in     vl_logic_vector;
        d116            : in     vl_logic_vector;
        d117            : in     vl_logic_vector;
        d118            : in     vl_logic_vector;
        d119            : in     vl_logic_vector;
        d120            : in     vl_logic_vector;
        d121            : in     vl_logic_vector;
        d122            : in     vl_logic_vector;
        d123            : in     vl_logic_vector;
        d124            : in     vl_logic_vector;
        d125            : in     vl_logic_vector;
        d126            : in     vl_logic_vector;
        d127            : in     vl_logic_vector;
        d128            : in     vl_logic_vector;
        d129            : in     vl_logic_vector;
        d130            : in     vl_logic_vector;
        d131            : in     vl_logic_vector;
        d132            : in     vl_logic_vector;
        d133            : in     vl_logic_vector;
        d134            : in     vl_logic_vector;
        d135            : in     vl_logic_vector;
        d136            : in     vl_logic_vector;
        d137            : in     vl_logic_vector;
        d138            : in     vl_logic_vector;
        d139            : in     vl_logic_vector;
        d140            : in     vl_logic_vector;
        d141            : in     vl_logic_vector;
        d142            : in     vl_logic_vector;
        d143            : in     vl_logic_vector;
        d144            : in     vl_logic_vector;
        d145            : in     vl_logic_vector;
        d146            : in     vl_logic_vector;
        d147            : in     vl_logic_vector;
        d148            : in     vl_logic_vector;
        d149            : in     vl_logic_vector;
        d150            : in     vl_logic_vector;
        d151            : in     vl_logic_vector;
        d152            : in     vl_logic_vector;
        d153            : in     vl_logic_vector;
        d154            : in     vl_logic_vector;
        d155            : in     vl_logic_vector;
        d156            : in     vl_logic_vector;
        d157            : in     vl_logic_vector;
        d158            : in     vl_logic_vector;
        d159            : in     vl_logic_vector;
        d160            : in     vl_logic_vector;
        d161            : in     vl_logic_vector;
        d162            : in     vl_logic_vector;
        d163            : in     vl_logic_vector;
        d164            : in     vl_logic_vector;
        d165            : in     vl_logic_vector;
        d166            : in     vl_logic_vector;
        d167            : in     vl_logic_vector;
        d168            : in     vl_logic_vector;
        d169            : in     vl_logic_vector;
        d170            : in     vl_logic_vector;
        d171            : in     vl_logic_vector;
        d172            : in     vl_logic_vector;
        d173            : in     vl_logic_vector;
        d174            : in     vl_logic_vector;
        d175            : in     vl_logic_vector;
        d176            : in     vl_logic_vector;
        d177            : in     vl_logic_vector;
        d178            : in     vl_logic_vector;
        d179            : in     vl_logic_vector;
        d180            : in     vl_logic_vector;
        d181            : in     vl_logic_vector;
        d182            : in     vl_logic_vector;
        d183            : in     vl_logic_vector;
        d184            : in     vl_logic_vector;
        d185            : in     vl_logic_vector;
        d186            : in     vl_logic_vector;
        d187            : in     vl_logic_vector;
        d188            : in     vl_logic_vector;
        d189            : in     vl_logic_vector;
        d190            : in     vl_logic_vector;
        d191            : in     vl_logic_vector;
        d192            : in     vl_logic_vector;
        d193            : in     vl_logic_vector;
        d194            : in     vl_logic_vector;
        d195            : in     vl_logic_vector;
        d196            : in     vl_logic_vector;
        d197            : in     vl_logic_vector;
        d198            : in     vl_logic_vector;
        d199            : in     vl_logic_vector;
        d200            : in     vl_logic_vector;
        d201            : in     vl_logic_vector;
        d202            : in     vl_logic_vector;
        d203            : in     vl_logic_vector;
        d204            : in     vl_logic_vector;
        d205            : in     vl_logic_vector;
        d206            : in     vl_logic_vector;
        d207            : in     vl_logic_vector;
        d208            : in     vl_logic_vector;
        d209            : in     vl_logic_vector;
        d210            : in     vl_logic_vector;
        d211            : in     vl_logic_vector;
        d212            : in     vl_logic_vector;
        d213            : in     vl_logic_vector;
        d214            : in     vl_logic_vector;
        d215            : in     vl_logic_vector;
        d216            : in     vl_logic_vector;
        d217            : in     vl_logic_vector;
        d218            : in     vl_logic_vector;
        d219            : in     vl_logic_vector;
        d220            : in     vl_logic_vector;
        d221            : in     vl_logic_vector;
        d222            : in     vl_logic_vector;
        d223            : in     vl_logic_vector;
        d224            : in     vl_logic_vector;
        d225            : in     vl_logic_vector;
        d226            : in     vl_logic_vector;
        d227            : in     vl_logic_vector;
        d228            : in     vl_logic_vector;
        d229            : in     vl_logic_vector;
        d230            : in     vl_logic_vector;
        d231            : in     vl_logic_vector;
        d232            : in     vl_logic_vector;
        d233            : in     vl_logic_vector;
        d234            : in     vl_logic_vector;
        d235            : in     vl_logic_vector;
        d236            : in     vl_logic_vector;
        d237            : in     vl_logic_vector;
        d238            : in     vl_logic_vector;
        d239            : in     vl_logic_vector;
        d240            : in     vl_logic_vector;
        d241            : in     vl_logic_vector;
        d242            : in     vl_logic_vector;
        d243            : in     vl_logic_vector;
        d244            : in     vl_logic_vector;
        d245            : in     vl_logic_vector;
        d246            : in     vl_logic_vector;
        d247            : in     vl_logic_vector;
        d248            : in     vl_logic_vector;
        d249            : in     vl_logic_vector;
        d250            : in     vl_logic_vector;
        d251            : in     vl_logic_vector;
        d252            : in     vl_logic_vector;
        d253            : in     vl_logic_vector;
        d254            : in     vl_logic_vector;
        d255            : in     vl_logic_vector;
        s               : in     vl_logic_vector(7 downto 0);
        y               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of WIDTH : constant is 1;
end mux255;
